`define OR or #20

module ALUor 
(
    output[31:0] oroutput,
    input[31:0] A,
    input[31:0] B
);

`OR orgate0(oroutput[0], A[0], B[0]);
`OR orgate1(oroutput[1], A[1], B[1]);
`OR orgate2(oroutput[2], A[2], B[2]);
`OR orgate3(oroutput[3], A[3], B[3]);
`OR orgate4(oroutput[4], A[4], B[4]);
`OR orgate5(oroutput[5], A[5], B[5]);
`OR orgate6(oroutput[6], A[6], B[6]);
`OR orgate7(oroutput[7], A[7], B[7]);
`OR orgate8(oroutput[8], A[8], B[8]);
`OR orgate9(oroutput[9], A[9], B[9]);
`OR orgate10(oroutput[10], A[10], B[10]);
`OR orgate11(oroutput[11], A[11], B[11]);
`OR orgate12(oroutput[12], A[12], B[12]);
`OR orgate13(oroutput[13], A[13], B[13]);
`OR orgate14(oroutput[14], A[14], B[14]);
`OR orgate15(oroutput[15], A[15], B[15]);
`OR orgate16(oroutput[16], A[16], B[16]);
`OR orgate17(oroutput[17], A[17], B[17]);
`OR orgate18(oroutput[18], A[18], B[18]);
`OR orgate19(oroutput[19], A[19], B[19]);
`OR orgate20(oroutput[20], A[20], B[20]);
`OR orgate21(oroutput[21], A[21], B[21]);
`OR orgate22(oroutput[22], A[22], B[22]);
`OR orgate23(oroutput[23], A[23], B[23]);
`OR orgate24(oroutput[24], A[24], B[24]);
`OR orgate25(oroutput[25], A[25], B[25]);
`OR orgate26(oroutput[26], A[26], B[26]);
`OR orgate27(oroutput[27], A[27], B[27]);
`OR orgate28(oroutput[28], A[28], B[28]);
`OR orgate29(oroutput[29], A[29], B[29]);
`OR orgate30(oroutput[30], A[30], B[30]);
`OR orgate31(oroutput[31], A[31], B[31]);

endmodule

