`define AND and #20

module ALUand
(
    output[31:0] andoutput,
    input[31:0] A,
    input[31:0] B
);

`AND andgate0(andoutput[0], A[0], B[0]);
`AND andgate1(andoutput[1], A[1], B[1]);
`AND andgate2(andoutput[2], A[2], B[2]);
`AND andgate3(andoutput[3], A[3], B[3]);
`AND andgate4(andoutput[4], A[4], B[4]);
`AND andgate5(andoutput[5], A[5], B[5]);
`AND andgate6(andoutput[6], A[6], B[6]);
`AND andgate7(andoutput[7], A[7], B[7]);
`AND andgate8(andoutput[8], A[8], B[8]);
`AND andgate9(andoutput[9], A[9], B[9]);
`AND andgate10(andoutput[10], A[10], B[10]);
`AND andgate11(andoutput[11], A[11], B[11]);
`AND andgate12(andoutput[12], A[12], B[12]);
`AND andgate13(andoutput[13], A[13], B[13]);
`AND andgate14(andoutput[14], A[14], B[14]);
`AND andgate15(andoutput[15], A[15], B[15]);
`AND andgate16(andoutput[16], A[16], B[16]);
`AND andgate17(andoutput[17], A[17], B[17]);
`AND andgate18(andoutput[18], A[18], B[18]);
`AND andgate19(andoutput[19], A[19], B[19]);
`AND andgate20(andoutput[20], A[20], B[20]);
`AND andgate21(andoutput[21], A[21], B[21]);
`AND andgate22(andoutput[22], A[22], B[22]);
`AND andgate23(andoutput[23], A[23], B[23]);
`AND andgate24(andoutput[24], A[24], B[24]);
`AND andgate25(andoutput[25], A[25], B[25]);
`AND andgate26(andoutput[26], A[26], B[26]);
`AND andgate27(andoutput[27], A[27], B[27]);
`AND andgate28(andoutput[28], A[28], B[28]);
`AND andgate29(andoutput[29], A[29], B[29]);
`AND andgate30(andoutput[30], A[30], B[30]);
`AND andgate31(andoutput[31], A[31], B[31]);

endmodule
